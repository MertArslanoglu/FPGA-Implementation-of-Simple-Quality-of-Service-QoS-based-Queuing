library verilog;
use verilog.vl_types.all;
entity proje_vlg_vec_tst is
end proje_vlg_vec_tst;
